library verilog;
use verilog.vl_types.all;
entity SYNC_COUNTER_vlg_vec_tst is
end SYNC_COUNTER_vlg_vec_tst;
