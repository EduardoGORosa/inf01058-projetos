library verilog;
use verilog.vl_types.all;
entity CODER_vlg_vec_tst is
end CODER_vlg_vec_tst;
