library verilog;
use verilog.vl_types.all;
entity Mux8bits21_vlg_vec_tst is
end Mux8bits21_vlg_vec_tst;
