library verilog;
use verilog.vl_types.all;
entity comp_igual_vlg_vec_tst is
end comp_igual_vlg_vec_tst;
