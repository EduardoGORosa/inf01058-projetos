library verilog;
use verilog.vl_types.all;
entity TrafficLights_vlg_vec_tst is
end TrafficLights_vlg_vec_tst;
