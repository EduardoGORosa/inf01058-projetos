library verilog;
use verilog.vl_types.all;
entity mux4bits21_vlg_vec_tst is
end mux4bits21_vlg_vec_tst;
