library verilog;
use verilog.vl_types.all;
entity ULA_DISPLAY_vlg_sample_tst is
    port(
        a               : in     vl_logic_vector(3 downto 0);
        b               : in     vl_logic_vector(3 downto 0);
        s               : in     vl_logic_vector(1 downto 0);
        sampler_tx      : out    vl_logic
    );
end ULA_DISPLAY_vlg_sample_tst;
