library verilog;
use verilog.vl_types.all;
entity DECODER_vlg_vec_tst is
end DECODER_vlg_vec_tst;
