library verilog;
use verilog.vl_types.all;
entity ULA_DISPLAY_vlg_vec_tst is
end ULA_DISPLAY_vlg_vec_tst;
