library verilog;
use verilog.vl_types.all;
entity MUX2_1_8_vlg_vec_tst is
end MUX2_1_8_vlg_vec_tst;
